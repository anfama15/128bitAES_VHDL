library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity subword is
 Port (
        i_state : in  std_logic_vector(31 downto 0);
        o_state : out std_logic_vector(31 downto 0);
        rot_check : out std_logic_vector(31 downto 0)
    );
end subword;

architecture Behavioral of subword is
    component RotWord is port(
           key_in   :   IN  std_logic_vector    (31 downto 0);
           data_out :   OUT std_logic_vector    (31 downto 0)
    );
    end component;
signal rot_in :  std_logic_vector (31 downto 0);
signal rot_out :  std_logic_vector (31 downto 0);
 function SBox(i_byte: std_logic_vector(7 downto 0)) return std_logic_vector is
        variable sbox_val: std_logic_vector(7 downto 0);
    begin

    
        case i_byte is
            when x"00" => sbox_val := x"63";
            when x"01" => sbox_val := x"7c";
            when x"02" => sbox_val := x"77";
            when x"03" => sbox_val := x"7b";
            when x"04" => sbox_val := x"f2";
            when x"05" => sbox_val := x"6b";
            when x"06" => sbox_val := x"6f";
            when x"07" => sbox_val := x"c5";
            when x"08" => sbox_val := x"30";
            when x"09" => sbox_val := x"01";
            when x"0a" => sbox_val := x"67";
            when x"0b" => sbox_val := x"2b";
            when x"0c" => sbox_val := x"fe";
            when x"0d" => sbox_val := x"d7";
            when x"0e" => sbox_val := x"ab";
            when x"0f" => sbox_val := x"76";
            when x"10" => sbox_val := x"ca";
            when x"11" => sbox_val := x"82";
            when x"12" => sbox_val := x"c9";
            when x"13" => sbox_val := x"7d";
            when x"14" => sbox_val := x"fa";
            when x"15" => sbox_val := x"59";
            when x"16" => sbox_val := x"47";
            when x"17" => sbox_val := x"f0";
            when x"18" => sbox_val := x"ad";
            when x"19" => sbox_val := x"d4";
            when x"1a" => sbox_val := x"a2";
            when x"1b" => sbox_val := x"af";
            when x"1c" => sbox_val := x"9c";
            when x"1d" => sbox_val := x"a4";
            when x"1e" => sbox_val := x"72";
            when x"1f" => sbox_val := x"c0";
            when x"20" => sbox_val := x"b7";
            when x"21" => sbox_val := x"fd";
            when x"22" => sbox_val := x"93";
            when x"23" => sbox_val := x"26";
            when x"24" => sbox_val := x"36";
            when x"25" => sbox_val := x"3f";
            when x"26" => sbox_val := x"f7";
            when x"27" => sbox_val := x"cc";
            when x"28" => sbox_val := x"34";
            when x"29" => sbox_val := x"a5";
            when x"2a" => sbox_val := x"e5";
            when x"2b" => sbox_val := x"f1";
            when x"2c" => sbox_val := x"71";
            when x"2d" => sbox_val := x"d8";
            when x"2e" => sbox_val := x"31";
            when x"2f" => sbox_val := x"15";
            when x"30" => sbox_val := x"04";
            when x"31" => sbox_val := x"c7";
            when x"32" => sbox_val := x"23";
            when x"33" => sbox_val := x"c3";
            when x"34" => sbox_val := x"18";
            when x"35" => sbox_val := x"96";
            when x"36" => sbox_val := x"05";
            when x"37" => sbox_val := x"9a";
            when x"38" => sbox_val := x"07";
            when x"39" => sbox_val := x"12";
            when x"3a" => sbox_val := x"80";
            when x"3b" => sbox_val := x"e2";
            when x"3c" => sbox_val := x"eb";
            when x"3d" => sbox_val := x"27";
            when x"3e" => sbox_val := x"b2";
            when x"3f" => sbox_val := x"75";
            when x"40" => sbox_val := x"09";
            when x"41" => sbox_val := x"83";
            when x"42" => sbox_val := x"2c";
            when x"43" => sbox_val := x"1a";
            when x"44" => sbox_val := x"1b";
            when x"45" => sbox_val := x"6e";
            when x"46" => sbox_val := x"5a";
            when x"47" => sbox_val := x"a0";
            when x"48" => sbox_val := x"52";
            when x"49" => sbox_val := x"3b";
            when x"4a" => sbox_val := x"d6";
            when x"4b" => sbox_val := x"b3";
            when x"4c" => sbox_val := x"29";
            when x"4d" => sbox_val := x"e3";
            when x"4e" => sbox_val := x"2f";
            when x"4f" => sbox_val := x"84";
            when x"50" => sbox_val := x"53";
            when x"51" => sbox_val := x"d1";
            when x"52" => sbox_val := x"00";
            when x"53" => sbox_val := x"ed";
            when x"54" => sbox_val := x"20";
            when x"55" => sbox_val := x"fc";
            when x"56" => sbox_val := x"b1";
            when x"57" => sbox_val := x"5b";
            when x"58" => sbox_val := x"6a";
            when x"59" => sbox_val := x"cb";
            when x"5a" => sbox_val := x"be";
            when x"5b" => sbox_val := x"39";
            when x"5c" => sbox_val := x"4a";
            when x"5d" => sbox_val := x"4c";
            when x"5e" => sbox_val := x"58";
            when x"5f" => sbox_val := x"cf";
            when x"60" => sbox_val := x"d0";
            when x"61" => sbox_val := x"ef";
            when x"62" => sbox_val := x"aa";
            when x"63" => sbox_val := x"fb";
            when x"64" => sbox_val := x"43";
            when x"65" => sbox_val := x"4d";
            when x"66" => sbox_val := x"33";
            when x"67" => sbox_val := x"85";
            when x"68" => sbox_val := x"45";
            when x"69" => sbox_val := x"f9";
            when x"6a" => sbox_val := x"02";
            when x"6b" => sbox_val := x"7f";
            when x"6c" => sbox_val := x"50";
            when x"6d" => sbox_val := x"3c";
            when x"6e" => sbox_val := x"9f";
            when x"6f" => sbox_val := x"a8";
            when x"70" => sbox_val := x"51";
            when x"71" => sbox_val := x"a3";
            when x"72" => sbox_val := x"40";
            when x"73" => sbox_val := x"8f";
            when x"74" => sbox_val := x"92";
            when x"75" => sbox_val := x"9d";
            when x"76" => sbox_val := x"38";
            when x"77" => sbox_val := x"f5";
            when x"78" => sbox_val := x"bc";
            when x"79" => sbox_val := x"b6";
            when x"7a" => sbox_val := x"da";
            when x"7b" => sbox_val := x"21";
            when x"7c" => sbox_val := x"10";
            when x"7d" => sbox_val := x"ff";
            when x"7e" => sbox_val := x"f3";
            when x"7f" => sbox_val := x"d2";
            when x"80" => sbox_val := x"cd";
            when x"81" => sbox_val := x"0c";
            when x"82" => sbox_val := x"13";
            when x"83" => sbox_val := x"ec";
            when x"84" => sbox_val := x"5f";
            when x"85" => sbox_val := x"97";
            when x"86" => sbox_val := x"44";
            when x"87" => sbox_val := x"17";
            when x"88" => sbox_val := x"c4";
            when x"89" => sbox_val := x"a7";
            when x"8a" => sbox_val := x"7e";
            when x"8b" => sbox_val := x"3d";
            when x"8c" => sbox_val := x"64";
            when x"8d" => sbox_val := x"5d";
            when x"8e" => sbox_val := x"19";
            when x"8f" => sbox_val := x"73";
            when x"90" => sbox_val := x"60";
            when x"91" => sbox_val := x"81";
            when x"92" => sbox_val := x"4f";
            when x"93" => sbox_val := x"dc";
            when x"94" => sbox_val := x"22";
            when x"95" => sbox_val := x"2a";
            when x"96" => sbox_val := x"90";
            when x"97" => sbox_val := x"88";
            when x"98" => sbox_val := x"46";
            when x"99" => sbox_val := x"ee";
            when x"9a" => sbox_val := x"b8";
            when x"9b" => sbox_val := x"14";
            when x"9c" => sbox_val := x"de";
            when x"9d" => sbox_val := x"5e";
            when x"9e" => sbox_val := x"0b";
            when x"9f" => sbox_val := x"db";
            when x"a0" => sbox_val := x"e0";
            when x"a1" => sbox_val := x"32";
            when x"a2" => sbox_val := x"3a";
            when x"a3" => sbox_val := x"0a";
            when x"a4" => sbox_val := x"49";
            when x"a5" => sbox_val := x"06";
            when x"a6" => sbox_val := x"24";
            when x"a7" => sbox_val := x"5c";
            when x"a8" => sbox_val := x"c2";
            when x"a9" => sbox_val := x"d3";
            when x"aa" => sbox_val := x"ac";
            when x"ab" => sbox_val := x"62";
            when x"ac" => sbox_val := x"91";
            when x"ad" => sbox_val := x"95";
            when x"ae" => sbox_val := x"e4";
            when x"af" => sbox_val := x"79";
            when x"b0" => sbox_val := x"e7";
            when x"b1" => sbox_val := x"c8";
            when x"b2" => sbox_val := x"37";
            when x"b3" => sbox_val := x"6d";
            when x"b4" => sbox_val := x"8d";
            when x"b5" => sbox_val := x"d5";
            when x"b6" => sbox_val := x"4e";
            when x"b7" => sbox_val := x"a9";
            when x"b8" => sbox_val := x"6c";
            when x"b9" => sbox_val := x"56";
            when x"ba" => sbox_val := x"f4";
            when x"bb" => sbox_val := x"ea";
            when x"bc" => sbox_val := x"65";
            when x"bd" => sbox_val := x"7a";
            when x"be" => sbox_val := x"ae";
            when x"bf" => sbox_val := x"08";
            when x"c0" => sbox_val := x"ba";
            when x"c1" => sbox_val := x"78";
            when x"c2" => sbox_val := x"25";
            when x"c3" => sbox_val := x"2e";
            when x"c4" => sbox_val := x"1c";
            when x"c5" => sbox_val := x"a6";
            when x"c6" => sbox_val := x"b4";
            when x"c7" => sbox_val := x"c6";
            when x"c8" => sbox_val := x"e8";
            when x"c9" => sbox_val := x"dd";
            when x"ca" => sbox_val := x"74";
            when x"cb" => sbox_val := x"1f";
            when x"cc" => sbox_val := x"4b";
            when x"cd" => sbox_val := x"bd";
            when x"ce" => sbox_val := x"8b";
            when x"cf" => sbox_val := x"8a";
            when x"d0" => sbox_val := x"70";
            when x"d1" => sbox_val := x"3e";
            when x"d2" => sbox_val := x"b5";
            when x"d3" => sbox_val := x"66";
            when x"d4" => sbox_val := x"48";
            when x"d5" => sbox_val := x"03";
            when x"d6" => sbox_val := x"f6";
            when x"d7" => sbox_val := x"0e";
            when x"d8" => sbox_val := x"61";
            when x"d9" => sbox_val := x"35";
            when x"da" => sbox_val := x"57";
            when x"db" => sbox_val := x"b9";
            when x"dc" => sbox_val := x"86";
            when x"dd" => sbox_val := x"c1";
            when x"de" => sbox_val := x"1d";
            when x"df" => sbox_val := x"9e";
            when x"e0" => sbox_val := x"e1";
            when x"e1" => sbox_val := x"f8";
            when x"e2" => sbox_val := x"98";
            when x"e3" => sbox_val := x"11";
            when x"e4" => sbox_val := x"69";
            when x"e5" => sbox_val := x"d9";
            when x"e6" => sbox_val := x"8e";
            when x"e7" => sbox_val := x"94";
            when x"e8" => sbox_val := x"9b";
            when x"e9" => sbox_val := x"1e";
            when x"ea" => sbox_val := x"87";
            when x"eb" => sbox_val := x"e9";
            when x"ec" => sbox_val := x"ce";
            when x"ed" => sbox_val := x"55";
            when x"ee" => sbox_val := x"28";
            when x"ef" => sbox_val := x"df";
            when x"f0" => sbox_val := x"8c";
            when x"f1" => sbox_val := x"a1";
            when x"f2" => sbox_val := x"89";
            when x"f3" => sbox_val := x"0d";
            when x"f4" => sbox_val := x"bf";
            when x"f5" => sbox_val := x"e6";
            when x"f6" => sbox_val := x"42";
            when x"f7" => sbox_val := x"68";
            when x"f8" => sbox_val := x"41";
            when x"f9" => sbox_val := x"99";
            when x"fa" => sbox_val := x"2d";
            when x"fb" => sbox_val := x"0f";
            when x"fc" => sbox_val := x"b0";
            when x"fd" => sbox_val := x"54";
            when x"fe" => sbox_val := x"bb";
            when x"ff" => sbox_val := x"16";
            when others => sbox_val := (others => '0');
        end case;
        return sbox_val;
    end function;
signal temp1 : std_logic_vector(31 downto 0);
signal temp2 : std_logic_vector(31 downto 0);

begin

    R1 : RotWord Port map (
    key_in   => i_state,
    data_out => temp1
);
rot_check <= temp1;

-- i =0*8+7= 7
--0=7 downto 0;
--1=15 downto 8  ;
--(i*8+7 downto i*8);
    process(temp1)
        variable temp_state: std_logic_vector(31 downto 0);
        variable byte_in, byte_out: std_logic_vector(7 downto 0);
    begin
        for i in 0 to 3 loop
            byte_in := temp1(i*8+7 downto i*8);
            byte_out := SBox(byte_in);
            temp_state(i*8+7 downto i*8) := byte_out;
        end loop;
        o_state <= temp_state;
    end process;
end Behavioral;



